/*
 * file: tc_pkg.sv
 *
 */

package tb_pkg;
  
  const time CLK_PERIOD_HALF = 5ns;


endpackage