/*
 * file: tc_pkg.sv
 *
 */

package tb_pkg;
  
  const time CLK_PERIOD = 20ns;
  


endpackage