/*
 * file: logIP_ifs.sv
 *
 */

//
// Interface to control xon/xoff flow control
// of uart tx unit
//
interface FlowCtr;
  logic xon;
  logic xoff;
  logic stb;
  modport Master (output xon, output xoff, output stb);
  modport Slave (input xon, input xoff, input stb);
endinterface : FlowCtr




