/*
 * file: uart8.svh
 * usage: 
 * 
 */

`ifndef H_UART8
`define H_UART8

typedef byte uart_item_t;
typedef mailbox #(uart_item_t) mxb_uart_t;

`endif