/*
 * file: tc_pkg.sv
 *
 */
`timescale 1ns/1ps
package tb_pkg;
  
  const time CLK_PERIOD_HALF = 5;


endpackage