/*
 * file: logIP.sv
 * usage: Top level module for logIP.
 *
 */