
// TODO delete if not required for sim